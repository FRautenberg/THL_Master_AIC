** Profile: "lab3 optimzed-dc sweep"  [ c:\users\finn\documents\github\master-thl-aic\lab_3\pspice\lab3-cascode-comparisson-PSpiceFiles\lab3 optimzed\dc sweep.sim ] 

** Creating circuit file "dc sweep.cir" 
** WARNING: THIS AUTOMATICALLY GENERATED FILE MAY BE OVERWRITTEN BY SUBSEQUENT SIMULATIONS

*Libraries: 
* Profile Libraries :
* Local Libraries :
.LIB "../../../MovedFiles/tsmc_250nm.lib" 
* From [PSPICE NETLIST] section of C:\Users\Finn\AppData\Roaming\SPB_Data\cdssetup\OrCAD_PSpice\17.2.0\PSpice.ini file:
.lib "nomd.lib" 

*Analysis directives: 
.DC LIN V_VDCout 0 3 0.01 
.OPTIONS ADVCONV
.PROBE64 V(alias(*)) I(alias(*)) W(alias(*)) D(alias(*)) NOISE(alias(*)) 
.INC "..\lab3 optimzed.net" 


.END
